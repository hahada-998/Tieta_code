`include "rs35m2c16s_g5_define.vh"
`include "pwrseq_define.vh"

parameter PEAVEY_SUPPORT = 1'b1;  //comment1,ph configuration

/*

*/
endmodule